* D:\UM\YEAR 2\SEM 2\KIE2001\E1\E1_Simulation.sch

* Schematics Version 9.1 - Web Update 1
* Sun Apr 10 14:26:47 2022



** Analysis setup **
.ac DEC 200 100 23k
.tran 0ns 0.005 0 10u
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "E1_Simulation.net"
.INC "E1_Simulation.als"


.probe


.END
